-- f_pulse.vhd
